* C:\Users\SriRamajayam\eSim-Workspace\3bit_counter\3bit_counter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/09/22 05:44:26

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ vinisha_3bit_counter		
Q2  clk Net-_C1-Pad2_ GND eSim_NPN		
Q1  GND Net-_C2-Pad2_ Net-_C1-Pad1_ eSim_NPN		
R1  Net-_R1-Pad1_ Net-_C1-Pad1_ 1k		
R4  Net-_R1-Pad1_ clk 1k		
R2  Net-_R1-Pad1_ Net-_C1-Pad2_ 100k		
R3  Net-_R1-Pad1_ Net-_C2-Pad2_ 100k		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 7.24u		
C2  clk Net-_C2-Pad2_ 7.24u		
v1  Net-_R1-Pad1_ GND 5		
U4  clk rst Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_2		
U2  clk plot_v1		
U3  rst plot_v1		
v2  rst GND pulse		
U5  Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ out2 out1 out0 dac_bridge_3		
U6  out2 plot_v1		
U7  out1 plot_v1		
U8  out0 plot_v1		

.end
